//Subject:      CO project 2 - Shift_Left_Two_32
//--------------------------------------------------------------------------------
//Version:     1
//--------------------------------------------------------------------------------
//Description: 
//--------------------------------------------------------------------------------

module Shift_Left_Two_32(
    data_i,
    data_o
);

//I/O ports                    
input [32-1:0] data_i;
output [32-1:0] data_o;

//shift left 2
assign data_o = data_i << 2;


endmodule

/*
module stimulus;

reg[32-1: 0] in;
wire[32-1: 0] out;

Shift_Left_Two_32 sl2(in, out);

initial
begin
	in = 31;
	#1 $display("%b %b", in, out);
	

	in = 16;
	#1 $display("%b %b", in, out);
end

endmodule
*/
